`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:46:23 10/21/2022 
// Design Name: 
// Module Name:    ALU_unit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
/* 
    * Assignment - 6
    * Problem - 3
    * Semester - 5 (Autumn)
    * Group - 56
    * Group members - Utsav Mehta (20CS10069) and Vibhu (20CS10072)
*/



// ALU module to compute the result and flags based on ALUop and ALUsel
module ALU_unit (
    input signed [31:0] a, 
    input signed [31:0] b, 
    input ALUsel, 
    input [4:0] ALUop, 
    output reg carry, 
    output reg zero, 
    output reg sign, 
    output reg [31:0] result
);

    // Stores carry generated by adder1
    wire temp_carry;

    // Stores 32-bit output of not, adder1, shifter, and, xor, mux1, mux2 respectively from left to right.
    wire [31:0] out_not, out_adder, out_shifter, out_and, out_xor, out_mux1, out_mux2, out_diff;

    mux_32_to_1 mux1 (.a(a), .b(32'd1), .select(ALUsel), .out(out_mux1));
    mux_32_to_1 mux2 (.a(b), .b(out_not), .select(ALUsel), .out(out_mux2));

    adder_32_bit adder (.a(out_mux1), .b(out_mux2), .c_in(1'b0), .c_out(temp_carry), .sum(out_adder));

    shifter shifter1 (.in(out_mux1), .shamt(out_mux2), .dir(ALUop[1]), .out(out_shifter), .arith_or_logic(ALUop[0]));

	 diff diff1(
			.a(a),
			.b(b),
			.out_diff(out_diff)
	 );

    assign out_not = ~b;
    assign out_and = out_mux1 & out_mux2;
    assign out_xor = out_mux1 ^ out_mux2;

    // result changes on change of any input signal
    always @(*) begin
        
        if(ALUop == 5'b00000)
            result = out_mux1;
				
        else if (ALUop == 5'b00001) begin
            carry = temp_carry;
            result = out_adder;
        end
		  
        else if (ALUop == 5'b00101)
            result = out_adder;
        
		  else if (ALUop == 5'b10101)
            result = out_adder;
        
		  else if (ALUop == 5'b00010)
            result = out_and;
        
		  else if (ALUop == 5'b00011)
            result = out_xor;
        
		  else if (ALUop[4:2] == 3'b010)
            result = out_shifter;
				
		  else if (ALUop == 5'b001111)
				result = out_diff;
        
		  else
            result = 32'd0;
				
    end

    // Flags change on change of result
    always @(result) begin

        if (!result)
            zero = 1'b1;
        
		  else 
            zero = 1'b0;

        sign = result[31];
    end
    
endmodule