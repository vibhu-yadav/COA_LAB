`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   11:41:05 11/09/2022
// Design Name:   miniRISC_wrapper
// Module Name:   /home/vibhu/KGPminiRISC/miniRISC_wrapper_test.v
// Project Name:  KGPminiRISC
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: miniRISC_wrapper
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module miniRISC_wrapper_test;

	// Outputs
	wire ;

	// Instantiate the Unit Under Test (UUT)
	miniRISC_wrapper uut (
		.()
	);

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

