`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:41:31 11/09/2022 
// Design Name: 
// Module Name:    diff_encoder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
/* 
    * Assignment - 6
    * Problem - 3
    * Semester - 5 (Autumn)
    * Group - 56
    * Group members - Utsav Mehta (20CS10069) and Vibhu (20CS10072)
*/

module encoder(in, out_diff);

    input [31:0] in;
    output reg [5:0] out_diff;

    always @(*) begin
        case (in)
            32'b00000000000000000000000000000000: out_diff = 6'b100000;
            32'b00000000000000000000000000000001: out_diff = 6'b000001;
            32'b00000000000000000000000000000010: out_diff = 6'b000010;
            32'b00000000000000000000000000000100: out_diff = 6'b000011;
            32'b00000000000000000000000000001000: out_diff = 6'b000100;
            32'b00000000000000000000000000010000: out_diff = 6'b000101;
            32'b00000000000000000000000000100000: out_diff = 6'b000110;
            32'b00000000000000000000000001000000: out_diff = 6'b000111;
            32'b00000000000000000000000010000000: out_diff = 6'b001000;
            32'b00000000000000000000000100000000: out_diff = 6'b001001;
            32'b00000000000000000000001000000000: out_diff = 6'b001010;
            32'b00000000000000000000010000000000: out_diff = 6'b001011;
            32'b00000000000000000000100000000000: out_diff = 6'b001100;
            32'b00000000000000000001000000000000: out_diff = 6'b001101;
            32'b00000000000000000010000000000000: out_diff = 6'b001110;
            32'b00000000000000000100000000000000: out_diff = 6'b001111;
            32'b00000000000000001000000000000000: out_diff = 6'b010000;
            32'b00000000000000010000000000000000: out_diff = 6'b010001;
            32'b00000000000000100000000000000000: out_diff = 6'b010010;
            32'b00000000000001000000000000000000: out_diff = 6'b010011;
            32'b00000000000010000000000000000000: out_diff = 6'b010100;
            32'b00000000000100000000000000000000: out_diff = 6'b010101;
            32'b00000000001000000000000000000000: out_diff = 6'b010110;
            32'b00000000010000000000000000000000: out_diff = 6'b010111;
            32'b00000000100000000000000000000000: out_diff = 6'b011000;
            32'b00000001000000000000000000000000: out_diff = 6'b011001;
            32'b00000010000000000000000000000000: out_diff = 6'b011010;
            32'b00000100000000000000000000000000: out_diff = 6'b011011;
            32'b00001000000000000000000000000000: out_diff = 6'b011100;
            32'b00010000000000000000000000000000: out_diff = 6'b011101;
            32'b00100000000000000000000000000000: out_diff = 6'b011110;
            32'b01000000000000000000000000000000: out_diff = 6'b011111;
            default: out_diff = 6'b011111;
        endcase
    end

endmodule