`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   14:26:27 08/26/2022
// Design Name:   full_adder
// Module Name:   C:/Users/Student/Asgn_3_Grp_56/tb_full_adder.v
// Project Name:  Asgn_3_Grp_56
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: full_adder
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

/* 

    * Assignment - 3
    * Problem - 1.b
    * Semester - 5 (Autumn)
    * Group - 56
    * Group members - Utsav Mehta (20CS10069) and Vibhu (20CS10072)

*/

module tb_full_adder;

    // Inputs and Outputs
    reg input_a, input_b, carry_in;
    wire sum, carry_out;

    // Module Instantiations (Unit Under Test)
    full_adder f_a(input_a, input_b, carry_in, sum, carry_out);

    initial begin
        
        $monitor ("a = %d, b = %d, carry_in = %d, sum = %d, carry_out = %d", input_a, input_b, carry_in, sum, carry_out);

        // Input values initialization
        input_a = 0;
		  input_b = 0;
		  carry_in = 0;
        #50;
        input_a = 0; 
		  input_b = 0;
		  carry_in = 1;
        #50;
        input_a = 0; 
		  input_b = 1;
		  carry_in = 0;
        #50;
        input_a = 0;
		  input_b = 1;
		  carry_in = 1;
        #50;
        input_a = 1;
		  input_b = 0;
		  carry_in = 0;
        #50;
        input_a = 1;
		  input_b = 0;
		  carry_in = 1;
        #50;
        input_a = 1;
		  input_b = 1;
		  carry_in = 0;
        #50;
        input_a = 1;
		  input_b = 1;
		  carry_in = 1;

    end

endmodule